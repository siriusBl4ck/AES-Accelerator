module aes(
    input [127:0] plaintxt_encrypt,
    output [127:0] ciphertxt_encrypt,
    input en_encrypt,
    output rdy_encrypt,
    input [127:0] ciphertxt_decrypt,
    output [127:0] plaintxt_decrypt,
    input en_decrypt,
    output rdy_decrypt
);
endmodule