module gf4_mult_t(input[3:0]x , input[3:0]y,output [3:0] out);

wire [6:0]c;
wire [6:0]d;
wire [6:0]out1;
assign c[0]=(x[0]&y[0]);
assign c[1]=(x[0]&y[1] ^ x[1]&y[0]);
assign c[2]=(x[0]&y[2] ^ x[1]&y[1] ^ x[2]&y[0]);
assign c[3]=(x[0]&y[3] ^ x[1]&y[2] ^ x[2]&y[1]  ^ x[3]&y[0]);
assign c[4]=(x[3]&y[1] ^ x[2]&y[2] ^ x[1]&y[3]);
assign c[5]=(x[3]&y[2] ^ x[2]&y[3]);
assign c[6]=(x[3]&y[3]);
assign out1[3]= (c[6]^c[3]) ;
assign out1[2]= (c[6] ^ c[5] ^  c[2] );
assign out1[1]= (c[5] ^ c[4] ^c[1] );
assign out1[0]= ((c[4]) ^c[0]);
assign d[0]=(out1[0]&1'b1);
assign d[1]=(out1[0]&1'b0^out1[1]&1'b1);
assign d[2]=(out1[0]&1'b0^out1[1]&1'b0^ out1[2]&1'b1);
assign d[3]=(out1[0]&1'b0^out1[1]&1'b0^ out1[2]&1'b0^out1[3]&1'b1);
assign d[4]=(out1[3]&1'b0^out1[2]&1'b0^ out1[1]&1'b0);
assign d[5]=(out1[3]&1'b0^out1[2]&1'b0);
assign d[6]=(out1[3]&1'b0);
assign out[3]= (d[6]^d[3]) ;
assign out[2]= (d[6] ^ d[5] ^ d[2] );
assign out[1]= (d[5] ^ d[4] ^d[1] );
assign out[0]= ((d[4]) ^d[0]);
endmodule